module IPS_tutorial (
    input signal,
    output LED
);

assing LED = ~signal;

endmodule


